module encoder4to2_tb;
    reg [3:0] in;
    wire [1:0] out;
    encoder4to2 uut(.in(in), .out(out));

    initial begin
        $monitor("in=%b => out=%b", in, out);
        in = 4'b0001; #10;
        in = 4'b0010; #10;
        in = 4'b0100; #10;
        in = 4'b1000; #10;
        $finish;
    end
endmodule



